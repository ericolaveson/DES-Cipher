//**********************************************************************************************************************
//* 
//* --------------------------------------------------------------------------------------------------------------------
//* 
//**********************************************************************************************************************
`ifndef _Definitions_v_
`define _Definitions_v_

typedef struct packed {
	logic [7:0] data;
} test_wire_s;

typedef test_wire_s t_wire;

`endif