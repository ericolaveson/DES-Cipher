/***********************************************************************************************************************
 * Eff Test Bench
 * ---------------------------------------------------------------------------------------------------------------------
 * This module will test the entire DES f function which folds the key into the cipher text and computes the DES
 * inverse.
 **********************************************************************************************************************/
`timescale 1ns / 1ps
`include "Definitions.sv"

module S_Boxes_tb #();

	logic clk; // clock signal
	
	// INITIALIZE - DES S_Box lines
	logic [47:0] s_wires_in;
	logic [3:0]  s_wires_out;
	
	// INITIALIZE - modules for testing
	S_Boxes  s_dut(s_wires_in, s_wires_out);
	
	
	// toggle the clock
	always begin
		#50ps  clk = 1;
		#50ps  clk = 0;
	end
	
	
	/*******************************************************************************************************************
	 *  _______ ______  _____ _______    _____ ______ ____  _    _ ______ _   _  _____ ______ 
	 * |__   __|  ____|/ ____|__   __|  / ____|  ____/ __ \| |  | |  ____| \ | |/ ____|  ____|
     *    | |  | |__  | (___    | |    | (___ | |__ | |  | | |  | | |__  |  \| | |    | |__   
     *    | |  |  __|  \___ \   | |     \___ \|  __|| |  | | |  | |  __| | . ` | |    |  __|  
     *    | |  | |____ ____) |  | |     ____) | |___| |__| | |__| | |____| |\  | |____| |____ 
     *    |_|  |______|_____/   |_|    |_____/|______\___\_\\____/|______|_| \_|\_____|______|
	 ******************************************************************************************************************/
	initial begin : test_S_Boxes
			clk        = 0;
			s_wires_in = 0;
		
		// TEST - set the input wires for test modules
		@(negedge clk);
		//                   000000000000000000000000000000000000000000000000
			s_wires_in = 48'b000000000000000000000000000000000000000010000000;
		
		repeat(20) @(negedge clk);
		
		$stop;
		
	end : test_S_Boxes
	
	
endmodule





















